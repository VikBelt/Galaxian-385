//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//                                                                       --
//    Fall 2014 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 7                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------

`include "game_params.sv"
import GAME_PARAMS::*;

module  color_mapper ( 
	input logic Clk, Reset, frame_clk, 
	input logic [7:0] keycode, 
	input [9:0] BallX, BallY, DrawX, DrawY, Ball_size,
	input [9:0] Alien1X, Alien1Y, Alien1S,
	input [9:0] Alien2X,Alien2Y,Alien2S,
	input [9:0] Alien3X,Alien3Y,Alien3S,
	input [9:0] Alien4X,Alien4Y,Alien4S,
	input [9:0] Alien5X,Alien5Y,Alien5S,
	input [9:0] Alien6X,Alien6Y,Alien6S,
	input [9:0] Alien7X,Alien7Y,Alien7S,
	input [9:0] Alien8X,Alien8Y,Alien8S,
	input [9:0] Alien9X,Alien9Y,Alien9S,
	input [9:0] Alien10X,Alien10Y,Alien10S,
	input [9:0] Alien11X,Alien11Y,Alien11S,
	input [9:0] Alien12X,Alien12Y,Alien12S,
	input [9:0] MissileX, MissileY, MissileS,
	input [9:0] Alien1MissileX, Alien1MissileY, Alien1MissileS,
	input [9:0] Alien2MissileX,Alien2MissileY,Alien2MissileS,
	input [9:0] Alien3MissileX,Alien3MissileY,Alien3MissileS,
	input [9:0] Alien4MissileX,Alien4MissileY,Alien4MissileS,
	input [9:0] Alien5MissileX,Alien5MissileY,Alien5MissileS,
	input [9:0] Alien6MissileX,Alien6MissileY,Alien6MissileS,
	input [9:0] Alien7MissileX,Alien7MissileY,Alien7MissileS,
	input [9:0] Alien8MissileX,Alien8MissileY,Alien8MissileS,
	input [9:0] Alien9MissileX,Alien9MissileY,Alien9MissileS,
	input [9:0] Alien10MissileX,Alien10MissileY,Alien10MissileS,
	input [9:0] Alien11MissileX,Alien11MissileY,Alien11MissileS,
	input [9:0] Alien12MissileX,Alien12MissileY,Alien12MissileS,
	input alien1_hit, 
	input alien2_hit, 
	input alien3_hit, 
	input alien4_hit, 
	input alien5_hit, 
	input alien6_hit, 
	input alien7_hit, 
	input alien8_hit, 
	input alien9_hit, 
	input alien10_hit, 
	input alien11_hit, 
	input alien12_hit,
	input missile_sight,
	input am1_sight,
	input am2_sight,
	input am3_sight,
	input am4_sight,
	input am5_sight,
	input am6_sight,
	input am7_sight,
	input am8_sight,
	input am9_sight,
	input am10_sight,
	input am11_sight,
	input am12_sight,
	input color_switch,
   output logic [7:0]  Red, Green, Blue 
);
    
	 /////////starfield generation/////////
	 //row one
	 logic star1_on, star2_on, star3_on, star4_on, star5_on, star6_on, star7_on, star8_on, star9_on, star10_on, star11_on, star12_on; //row one
	 int DistStar1X, DistStar1Y;
	 assign DistStar1X = DrawX - star_OneX;
	 assign DistStar1Y = DrawY - star_row_one;
	 
	 int DistStar2X, DistStar2Y;
	 assign DistStar2X = DrawX - star2_X;
	 assign DistStar2Y = DrawY - star_row_one;
	 
	 int DistStar3X, DistStar3Y;
	 assign DistStar3X = DrawX - star3_X;
	 assign DistStar3Y = DrawY - star_row_one;
	 
	 int DistStar4X, DistStar4Y;
	 assign DistStar4X = DrawX - star4_X;
	 assign DistStar4Y = DrawY - star_row_one;
	 
	 int DistStar5X, DistStar5Y;
	 assign DistStar5X = DrawX - star5_X;
	 assign DistStar5Y = DrawY - star_row_one;
	 
	 int DistStar6X, DistStar6Y;
	 assign DistStar6X = DrawX - star6_X;
	 assign DistStar6Y = DrawY - star_row_one;
	 
	 int DistStar7X, DistStar7Y;
	 assign DistStar7X = DrawX - star7_X;
	 assign DistStar7Y = DrawY - star_row_one;
	 
	 int DistStar8X, DistStar8Y;
	 assign DistStar8X = DrawX - star8_X;
	 assign DistStar8Y = DrawY - star_row_one;
	 
	 int DistStar9X, DistStar9Y;
	 assign DistStar9X = DrawX - star9_X;
	 assign DistStar9Y = DrawY - star_row_one;
	 
	 int DistStar10X, DistStar10Y;
	 assign DistStar10X = DrawX - star10_X;
	 assign DistStar10Y = DrawY - star_row_one;

	 int DistStar11X, DistStar11Y;
	 assign DistStar11X = DrawX - star11_X;
	 assign DistStar11Y = DrawY - star_row_one;
	 
	 int DistStar12X, DistStar12Y;
	 assign DistStar12X = DrawX - star12_X;
	 assign DistStar12Y = DrawY - star_row_one;
	 
	 //row two
	 logic star13_on, star14_on, star15_on, star16_on, star17_on, star18_on, star19_on, star20_on, star21_on, star22_on, star23_on, star24_on; //row two
	 int DistStar13X, DistStar13Y;
	 assign DistStar13X = DrawX - starB_OneX;
	 assign DistStar13Y = DrawY - star_row_two;
	 
	 int DistStar14X, DistStar14Y;
	 assign DistStar14X = DrawX - starB2_X;
	 assign DistStar14Y = DrawY - star_row_two;
	 
	 int DistStar15X, DistStar15Y;
	 assign DistStar15X = DrawX - starB3_X;
	 assign DistStar15Y = DrawY - star_row_two;
	 
	 int DistStar16X, DistStar16Y;
	 assign DistStar16X = DrawX - starB4_X;
	 assign DistStar16Y = DrawY - star_row_two;
	 
	 int DistStar17X, DistStar17Y;
	 assign DistStar17X = DrawX - starB5_X;
	 assign DistStar17Y = DrawY - star_row_two;
	 
	 int DistStar18X, DistStar18Y;
	 assign DistStar18X = DrawX - starB6_X;
	 assign DistStar18Y = DrawY - star_row_two;
	 
	 int DistStar19X, DistStar19Y;
	 assign DistStar19X = DrawX - starB7_X;
	 assign DistStar19Y = DrawY - star_row_two;
	 
	 int DistStar20X, DistStar20Y;
	 assign DistStar20X = DrawX - starB8_X;
	 assign DistStar20Y = DrawY - star_row_two;
	 
	 int DistStar21X, DistStar21Y;
	 assign DistStar21X = DrawX - starB9_X;
	 assign DistStar21Y = DrawY - star_row_two;
	 
	 int DistStar22X, DistStar22Y;
	 assign DistStar22X = DrawX - starB10_X;
	 assign DistStar22Y = DrawY - star_row_two;

	 int DistStar23X, DistStar23Y;
	 assign DistStar23X = DrawX - starB11_X;
	 assign DistStar23Y = DrawY - star_row_two;
	 
	 int DistStar24X, DistStar24Y;
	 assign DistStar24X = DrawX - starB12_X;
	 assign DistStar24Y = DrawY - star_row_two;
	 
	 //row three
	 logic star25_on, star26_on, star27_on, star28_on, star29_on, star30_on, star31_on, star32_on, star33_on, star34_on, star35_on, star36_on; //row three
	 int DistStar25X, DistStar25Y;
	 assign DistStar25X = DrawX - star_OneX;
	 assign DistStar25Y = DrawY - star_row_three;
	 
	 int DistStar26X, DistStar26Y;
	 assign DistStar26X = DrawX - star2_X;
	 assign DistStar26Y = DrawY - star_row_three;
	 
	 int DistStar27X, DistStar27Y;
	 assign DistStar27X = DrawX - star3_X;
	 assign DistStar27Y = DrawY - star_row_three;
	 
	 int DistStar28X, DistStar28Y;
	 assign DistStar28X = DrawX - star4_X;
	 assign DistStar28Y = DrawY - star_row_three;
	 
	 int DistStar29X, DistStar29Y;
	 assign DistStar29X = DrawX - star5_X;
	 assign DistStar29Y = DrawY - star_row_three;
	 
	 int DistStar30X, DistStar30Y;
	 assign DistStar30X = DrawX - star6_X;
	 assign DistStar30Y = DrawY - star_row_three;
	 
	 int DistStar31X, DistStar31Y;
	 assign DistStar31X = DrawX - star7_X;
	 assign DistStar31Y = DrawY - star_row_three;
	 
	 int DistStar32X, DistStar32Y;
	 assign DistStar32X = DrawX - star8_X;
	 assign DistStar32Y = DrawY - star_row_three;
	 
	 int DistStar33X, DistStar33Y;
	 assign DistStar33X = DrawX - star9_X;
	 assign DistStar33Y = DrawY - star_row_three;
	 
	 int DistStar34X, DistStar34Y;
	 assign DistStar34X = DrawX - star10_X;
	 assign DistStar34Y = DrawY - star_row_three;

	 int DistStar35X, DistStar35Y;
	 assign DistStar35X = DrawX - star11_X;
	 assign DistStar35Y = DrawY - star_row_three;
	 
	 int DistStar36X, DistStar36Y;
	 assign DistStar36X = DrawX - star12_X;
	 assign DistStar36Y = DrawY - star_row_three;
	 
    //row four
	 logic star37_on, star38_on, star39_on, star40_on, star41_on, star42_on, star43_on, star44_on, star45_on, star46_on, star47_on, star48_on; //row four
	 
	 int DistStar37X, DistStar37Y;
	 assign DistStar37X = DrawX - starB_OneX;
	 assign DistStar37Y = DrawY - star_row_four;
	 
	 int DistStar38X, DistStar38Y;
	 assign DistStar38X = DrawX - starB2_X;
	 assign DistStar38Y = DrawY - star_row_four;
	 
	 int DistStar39X, DistStar39Y;
	 assign DistStar39X = DrawX - starB3_X;
	 assign DistStar39Y = DrawY - star_row_four;
	 
	 int DistStar40X, DistStar40Y;
	 assign DistStar40X = DrawX - starB4_X;
	 assign DistStar40Y = DrawY - star_row_four;
	 
	 int DistStar41X, DistStar41Y;
	 assign DistStar41X = DrawX - starB5_X;
	 assign DistStar41Y = DrawY - star_row_four;
	 
	 int DistStar42X, DistStar42Y;
	 assign DistStar42X = DrawX - starB6_X;
	 assign DistStar42Y = DrawY - star_row_four;
	 
	 int DistStar43X, DistStar43Y;
	 assign DistStar43X = DrawX - starB7_X;
	 assign DistStar43Y = DrawY - star_row_four;
	 
	 int DistStar44X, DistStar44Y;
	 assign DistStar44X = DrawX - starB8_X;
	 assign DistStar44Y = DrawY - star_row_four;
	 
	 int DistStar45X, DistStar45Y;
	 assign DistStar45X = DrawX - starB9_X;
	 assign DistStar45Y = DrawY - star_row_four;
	 
	 int DistStar46X, DistStar46Y;
	 assign DistStar46X = DrawX - starB10_X;
	 assign DistStar46Y = DrawY - star_row_four;

	 int DistStar47X, DistStar47Y;
	 assign DistStar47X = DrawX - starB11_X;
	 assign DistStar47Y = DrawY - star_row_four;
	 
	 int DistStar48X, DistStar48Y;
	 assign DistStar48X = DrawX - starB12_X;
	 assign DistStar48Y = DrawY - star_row_four;

	 //row five
	 logic star49_on, star50_on, star51_on, star52_on, star53_on, star54_on, star55_on, star56_on, star57_on, star58_on, star59_on, star60_on; //row five
	 
	 int DistStar49X, DistStar49Y;
	 assign DistStar49X = DrawX - star_OneX;
	 assign DistStar49Y = DrawY - star_row_five;
	 
	 int DistStar50X, DistStar50Y;
	 assign DistStar50X = DrawX - star2_X;
	 assign DistStar50Y = DrawY - star_row_five;
	 
	 int DistStar51X, DistStar51Y;
	 assign DistStar51X = DrawX - star3_X;
	 assign DistStar51Y = DrawY - star_row_five;
	 
	 int DistStar52X, DistStar52Y;
	 assign DistStar52X = DrawX - star4_X;
	 assign DistStar52Y = DrawY - star_row_five;
	 
	 int DistStar53X, DistStar53Y;
	 assign DistStar53X = DrawX - star5_X;
	 assign DistStar53Y = DrawY - star_row_five;
	 
	 int DistStar54X, DistStar54Y;
	 assign DistStar54X = DrawX - star6_X;
	 assign DistStar54Y = DrawY - star_row_five;
	 
	 int DistStar55X, DistStar55Y;
	 assign DistStar55X = DrawX - star7_X;
	 assign DistStar55Y = DrawY - star_row_five;
	 
	 int DistStar56X, DistStar56Y;
	 assign DistStar56X = DrawX - star8_X;
	 assign DistStar56Y = DrawY - star_row_five;
	 
	 int DistStar57X, DistStar57Y;
	 assign DistStar57X = DrawX - star9_X;
	 assign DistStar57Y = DrawY - star_row_five;
	 
	 int DistStar58X, DistStar58Y;
	 assign DistStar58X = DrawX - star10_X;
	 assign DistStar58Y = DrawY - star_row_five;

	 int DistStar59X, DistStar59Y;
	 assign DistStar59X = DrawX - star11_X;
	 assign DistStar59Y = DrawY - star_row_five;
	 
	 int DistStar60X, DistStar60Y;
	 assign DistStar60X = DrawX - star12_X;
	 assign DistStar60Y = DrawY - star_row_five;

	 //row six
	 logic star61_on, star62_on, star63_on, star64_on, star65_on, star66_on, star67_on, star68_on, star69_on, star70_on, star71_on, star72_on; //row six
	 
	 int DistStar61X, DistStar61Y;
	 assign DistStar61X = DrawX - starB_OneX;
	 assign DistStar61Y = DrawY - star_row_six;
	 
	 int DistStar62X, DistStar62Y;
	 assign DistStar62X = DrawX - starB2_X;
	 assign DistStar62Y = DrawY - star_row_six;
	 
	 int DistStar63X, DistStar63Y;
	 assign DistStar63X = DrawX - starB3_X;
	 assign DistStar63Y = DrawY - star_row_six;
	 
	 int DistStar64X, DistStar64Y;
	 assign DistStar64X = DrawX - starB4_X;
	 assign DistStar64Y = DrawY - star_row_six;
	 
	 int DistStar65X, DistStar65Y;
	 assign DistStar65X = DrawX - starB5_X;
	 assign DistStar65Y = DrawY - star_row_six;
	 
	 int DistStar66X, DistStar66Y;
	 assign DistStar66X = DrawX - starB6_X;
	 assign DistStar66Y = DrawY - star_row_six;
	 
	 int DistStar67X, DistStar67Y;
	 assign DistStar67X = DrawX - starB7_X;
	 assign DistStar67Y = DrawY - star_row_six;
	 
	 int DistStar68X, DistStar68Y;
	 assign DistStar68X = DrawX - starB8_X;
	 assign DistStar68Y = DrawY - star_row_six;
	 
	 int DistStar69X, DistStar69Y;
	 assign DistStar69X = DrawX - starB9_X;
	 assign DistStar69Y = DrawY - star_row_six;
	 
	 int DistStar70X, DistStar70Y;
	 assign DistStar70X = DrawX - starB10_X;
	 assign DistStar70Y = DrawY - star_row_six;

	 int DistStar71X, DistStar71Y;
	 assign DistStar71X = DrawX - starB11_X;
	 assign DistStar71Y = DrawY - star_row_six;
	 
	 int DistStar72X, DistStar72Y;
	 assign DistStar72X = DrawX - starB12_X;
	 assign DistStar72Y = DrawY - star_row_six;

	 //row seven
	 logic star73_on, star74_on, star75_on, star76_on, star77_on, star78_on, star79_on, star80_on, star81_on, star82_on, star83_on, star84_on; //row seven
	 
	 int DistStar73X, DistStar73Y;
	 assign DistStar73X = DrawX - star_OneX;
	 assign DistStar73Y = DrawY - star_row_seven;
	 
	 int DistStar74X, DistStar74Y;
	 assign DistStar74X = DrawX - star2_X;
	 assign DistStar74Y = DrawY - star_row_seven;
	 
	 int DistStar75X, DistStar75Y;
	 assign DistStar75X = DrawX - star3_X;
	 assign DistStar75Y = DrawY - star_row_seven;
	 
	 int DistStar76X, DistStar76Y;
	 assign DistStar76X = DrawX - star4_X;
	 assign DistStar76Y = DrawY - star_row_seven;
	 
	 int DistStar77X, DistStar77Y;
	 assign DistStar77X = DrawX - star5_X;
	 assign DistStar77Y = DrawY - star_row_seven;
	 
	 int DistStar78X, DistStar78Y;
	 assign DistStar78X = DrawX - star6_X;
	 assign DistStar78Y = DrawY - star_row_seven;
	 
	 int DistStar79X, DistStar79Y;
	 assign DistStar79X = DrawX - star7_X;
	 assign DistStar79Y = DrawY - star_row_seven;
	 
	 int DistStar80X, DistStar80Y;
	 assign DistStar80X = DrawX - star8_X;
	 assign DistStar80Y = DrawY - star_row_seven;
	 
	 int DistStar81X, DistStar81Y;
	 assign DistStar81X = DrawX - star9_X;
	 assign DistStar81Y = DrawY - star_row_seven;
	 
	 int DistStar82X, DistStar82Y;
	 assign DistStar82X = DrawX - star10_X;
	 assign DistStar82Y = DrawY - star_row_seven;

	 int DistStar83X, DistStar83Y;
	 assign DistStar83X = DrawX - star11_X;
	 assign DistStar83Y = DrawY - star_row_seven;
	 
	 int DistStar84X, DistStar84Y;
	 assign DistStar84X = DrawX - star12_X;
	 assign DistStar84Y = DrawY - star_row_seven;

	 //row eight
	 logic star85_on, star86_on, star87_on, star88_on, star89_on, star90_on, star91_on, star92_on, star93_on, star94_on, star95_on, star96_on; //row eight
	 
	 int DistStar85X, DistStar85Y;
	 assign DistStar85X = DrawX - starB_OneX;
	 assign DistStar85Y = DrawY - star_row_eight;
	 
	 int DistStar86X, DistStar86Y;
	 assign DistStar86X = DrawX - starB2_X;
	 assign DistStar86Y = DrawY - star_row_eight;
	 
	 int DistStar87X, DistStar87Y;
	 assign DistStar87X = DrawX - starB3_X;
	 assign DistStar87Y = DrawY - star_row_eight;
	 
	 int DistStar88X, DistStar88Y;
	 assign DistStar88X = DrawX - starB4_X;
	 assign DistStar88Y = DrawY - star_row_eight;
	 
	 int DistStar89X, DistStar89Y;
	 assign DistStar89X = DrawX - starB5_X;
	 assign DistStar89Y = DrawY - star_row_eight;
	 
	 int DistStar90X, DistStar90Y;
	 assign DistStar90X = DrawX - starB6_X;
	 assign DistStar90Y = DrawY - star_row_eight;
	 
	 int DistStar91X, DistStar91Y;
	 assign DistStar91X = DrawX - starB7_X;
	 assign DistStar91Y = DrawY - star_row_eight;
	 
	 int DistStar92X, DistStar92Y;
	 assign DistStar92X = DrawX - starB8_X;
	 assign DistStar92Y = DrawY - star_row_eight;
	 
	 int DistStar93X, DistStar93Y;
	 assign DistStar93X = DrawX - starB9_X;
	 assign DistStar93Y = DrawY - star_row_eight;
	 
	 int DistStar94X, DistStar94Y;
	 assign DistStar94X = DrawX - starB10_X;
	 assign DistStar94Y = DrawY - star_row_eight;

	 int DistStar95X, DistStar95Y;
	 assign DistStar95X = DrawX - starB11_X;
	 assign DistStar95Y = DrawY - star_row_eight;
	 
	 int DistStar96X, DistStar96Y;
	 assign DistStar96X = DrawX - starB12_X;
	 assign DistStar96Y = DrawY - star_row_eight;

    //row nine
	 logic star97_on, star98_on, star99_on, star100_on, star101_on, star102_on, star103_on, star104_on, star105_on, star106_on, star107_on, star108_on; //row nine
	 int DistStar97X, DistStar97Y;
	 assign DistStar97X = DrawX - star_OneX;
	 assign DistStar97Y = DrawY - star_row_nine;
	 
	 int DistStar98X, DistStar98Y;
	 assign DistStar98X = DrawX - star2_X;
	 assign DistStar98Y = DrawY - star_row_nine;
	 
	 int DistStar99X, DistStar99Y;
	 assign DistStar99X = DrawX - star3_X;
	 assign DistStar99Y = DrawY - star_row_nine;
	 
	 int DistStar100X, DistStar100Y;
	 assign DistStar100X = DrawX - star4_X;
	 assign DistStar100Y = DrawY - star_row_nine;
	 
	 int DistStar101X, DistStar101Y;
	 assign DistStar101X = DrawX - star5_X;
	 assign DistStar101Y = DrawY - star_row_nine;
	 
	 int DistStar102X, DistStar102Y;
	 assign DistStar102X = DrawX - star6_X;
	 assign DistStar102Y = DrawY - star_row_nine;
	 
	 int DistStar103X, DistStar103Y;
	 assign DistStar103X = DrawX - star7_X;
	 assign DistStar103Y = DrawY - star_row_nine;
	 
	 int DistStar104X, DistStar104Y;
	 assign DistStar104X = DrawX - star8_X;
	 assign DistStar104Y = DrawY - star_row_nine;
	 
	 int DistStar105X, DistStar105Y;
	 assign DistStar105X = DrawX - star9_X;
	 assign DistStar105Y = DrawY - star_row_nine;
	 
	 int DistStar106X, DistStar106Y;
	 assign DistStar106X = DrawX - star10_X;
	 assign DistStar106Y = DrawY - star_row_nine;

	 int DistStar107X, DistStar107Y;
	 assign DistStar107X = DrawX - star11_X;
	 assign DistStar107Y = DrawY - star_row_nine;
	 
	 int DistStar108X, DistStar108Y;
	 assign DistStar108X = DrawX - star12_X;
	 assign DistStar108Y = DrawY - star_row_nine;

//	 //row ten
    logic star109_on, star110_on, star111_on, star112_on, star113_on, star114_on, star115_on, star116_on, star117_on, star118_on, star119_on, star120_on; //row ten
	 
	 int DistStar109X, DistStar109Y;
	 assign DistStar109X = DrawX - starB_OneX;
	 assign DistStar109Y = DrawY - star_row_ten;
	 
	 int DistStar110X, DistStar110Y;
	 assign DistStar110X = DrawX - starB2_X;
	 assign DistStar110Y = DrawY - star_row_ten;
	 
	 int DistStar111X, DistStar111Y;
	 assign DistStar111X = DrawX - starB3_X;
	 assign DistStar111Y = DrawY - star_row_ten;
	 
	 int DistStar112X, DistStar112Y;
	 assign DistStar112X = DrawX - starB4_X;
	 assign DistStar112Y = DrawY - star_row_ten;
	 
	 int DistStar113X, DistStar113Y;
	 assign DistStar113X = DrawX - starB5_X;
	 assign DistStar113Y = DrawY - star_row_ten;
	 
	 int DistStar114X, DistStar114Y;
	 assign DistStar114X = DrawX - starB6_X;
	 assign DistStar114Y = DrawY - star_row_ten;
	 
	 int DistStar115X, DistStar115Y;
	 assign DistStar115X = DrawX - starB7_X;
	 assign DistStar115Y = DrawY - star_row_ten;
	 
	 int DistStar116X, DistStar116Y;
	 assign DistStar116X = DrawX - starB8_X;
	 assign DistStar116Y = DrawY - star_row_ten;
	 
	 int DistStar117X, DistStar117Y;
	 assign DistStar117X = DrawX - starB9_X;
	 assign DistStar117Y = DrawY - star_row_ten;
	 
	 int DistStar118X, DistStar118Y;
	 assign DistStar118X = DrawX - starB10_X;
	 assign DistStar118Y = DrawY - star_row_ten;

	 int DistStar119X, DistStar119Y;
	 assign DistStar119X = DrawX - starB11_X;
	 assign DistStar119Y = DrawY - star_row_ten;
	 
	 int DistStar120X, DistStar120Y;
	 assign DistStar120X = DrawX - starB12_X;
	 assign DistStar120Y = DrawY - star_row_ten;
	 //////////end starfield///////////
		
		
	 //ball and sprite info
    logic ball_on;
	 logic [10:0] sprite_addr;
	 logic [7:0] sprite_data;

	 //declaring a new instance of the font_rom module (provided code)
	 font_rom(
		.addr(sprite_addr),
		.data(sprite_data)
	 );


	logic [18:0] ship_addr; 
	logic [23:0] dout;
	frameRAM ship_ram
	(
		.data_In(24'b0),
		.write_address(19'b0), 
		.read_address(ship_addr),
		.we(1'b0), 
		.Clk(Clk),
		.data_Out(dout)
	);
	
	logic [18:0] alien_addr; 
	logic [23:0] dout_1;
	alienRAM alien_ram
	(
		.data_In(24'b0),
		.write_address(19'b0), 
		.read_address(alien_addr),
		.we(1'b0), 
		.Clk(Clk),
		.data_Out(dout_1)
	);
	
	 logic missile_on;
	 logic alien1_on, alien2_on, alien3_on, alien4_on, alien5_on, alien6_on, alien7_on, alien8_on, alien9_on, alien10_on, alien11_on, alien12_on;
	 logic am1_on, am2_on, am3_on, am4_on, am5_on, am6_on, am7_on, am8_on, am9_on, am10_on, am11_on, am12_on;
	 
	 //Ball params
    int DistX, DistY, Size;
	 int DistAlien1X, DistAlien1Y, DistAlien2X, DistAlien2Y, DistAlien3X, DistAlien3Y, DistAlien4X, DistAlien4Y, DistAlien5X, DistAlien5Y, DistAlien6X, DistAlien6Y, DistAlien7X, DistAlien7Y;
	 int DistAlien8X, DistAlien8Y, DistAlien9X, DistAlien9Y, DistAlien10X, DistAlien10Y, DistAlien11X, DistAlien11Y, DistAlien12X, DistAlien12Y;
	 
	 assign DistAlien1X = DrawX - Alien1X; 
	 assign DistAlien1Y = DrawY - Alien1Y; 

	 assign DistAlien2X = DrawX - Alien2X; 
	 assign DistAlien2Y = DrawY - Alien2Y;
	 
	 assign DistAlien3X = DrawX - Alien3X; 
	 assign DistAlien3Y = DrawY - Alien3Y;
	 
	 assign DistAlien4X = DrawX - Alien4X; 
	 assign DistAlien4Y = DrawY - Alien4Y;
	 
	 assign DistAlien5X = DrawX - Alien5X; 
	 assign DistAlien5Y = DrawY - Alien5Y;
	 
	 assign DistAlien6X = DrawX - Alien6X; 
	 assign DistAlien6Y = DrawY - Alien6Y;
	 
	 assign DistAlien7X = DrawX - Alien7X; 
	 assign DistAlien7Y = DrawY - Alien7Y;
	 
	 assign DistAlien8X = DrawX - Alien8X; 
	 assign DistAlien8Y = DrawY - Alien8Y;
	 
	 assign DistAlien9X = DrawX - Alien9X; 
	 assign DistAlien9Y = DrawY - Alien9Y;
	 
	 assign DistAlien10X = DrawX - Alien10X; 
	 assign DistAlien10Y = DrawY - Alien10Y;
	 
	 assign DistAlien11X = DrawX - Alien11X; 
	 assign DistAlien11Y = DrawY - Alien11Y;
	 
	 assign DistAlien12X = DrawX - Alien12X; 
	 assign DistAlien12Y = DrawY - Alien12Y;
	 
	 assign DistX = DrawX - BallX;
    assign DistY = DrawY - BallY;
    assign Size = Ball_size;
	  
	 always_comb
	 //ship
	 begin:Ball_on_proj
		if (DrawX >= BallX && DrawX < BallX + Ball_size &&
			DrawY >= BallY && DrawY < BallY + Ball_size)
		begin
           ball_on = 1'b1;
			  alien1_on = 1'b0;
			  alien2_on = 1'b0;
			  alien3_on = 1'b0;
			  alien4_on = 1'b0;
			  alien5_on = 1'b0;
			  alien6_on = 1'b0;
			  alien7_on = 1'b0;
			  alien8_on = 1'b0;
		     alien9_on = 1'b0;
			  alien10_on = 1'b0;
			  alien11_on = 1'b0;
			  alien12_on = 1'b0;
			  missile_on = 1'b0;
			  am1_on = 1'b0;
			  am2_on = 1'b0;
			  am3_on = 1'b0;
			  am4_on = 1'b0;
			  am5_on = 1'b0;
			  am6_on = 1'b0;
			  am7_on = 1'b0;
			  am8_on = 1'b0;
		     am9_on = 1'b0;
			  am10_on = 1'b0;
			  am11_on = 1'b0;
			  am12_on = 1'b0;
			  sprite_addr = 10'b0;
			  star1_on = 1'b0;
			  star2_on = 1'b0;
			  star3_on = 1'b0;
			  star4_on = 1'b0;
			  star5_on = 1'b0;
			  star6_on = 1'b0;
			  star7_on = 1'b0;
			  star8_on = 1'b0;
			  star9_on = 1'b0;
			  star10_on = 1'b0;
			  star11_on = 1'b0;
			  star12_on = 1'b0;
			  star13_on = 1'b0;
			  star14_on = 1'b0;
			  star15_on = 1'b0;
			  star16_on = 1'b0;
			  star17_on = 1'b0;
			  star18_on = 1'b0;
			  star19_on = 1'b0;
			  star20_on = 1'b0;
			  star21_on = 1'b0;
			  star22_on = 1'b0;
			  star23_on = 1'b0;
			  star24_on = 1'b0;	
			  star25_on = 1'b0;
			  star26_on = 1'b0;
			  star27_on = 1'b0;
			  star28_on = 1'b0;
			  star29_on = 1'b0;
			  star30_on = 1'b0;
			  star31_on = 1'b0;
			  star32_on = 1'b0;
			  star33_on = 1'b0;
			  star34_on = 1'b0;
			  star35_on = 1'b0;
			  star36_on = 1'b0;
			  star37_on = 1'b0;
			  star38_on = 1'b0;
			  star39_on = 1'b0;
			  star40_on = 1'b0;
			  star41_on = 1'b0;
			  star42_on = 1'b0;
			  star43_on = 1'b0;
			  star44_on = 1'b0;
			  star45_on = 1'b0;
			  star46_on = 1'b0;
			  star47_on = 1'b0;
			  star48_on = 1'b0;
			  star49_on = 1'b0;
			  star50_on = 1'b0;
			  star51_on = 1'b0;
			  star52_on = 1'b0;
			  star53_on = 1'b0;
			  star54_on = 1'b0;
			  star55_on = 1'b0;
			  star56_on = 1'b0;
			  star57_on = 1'b0;
			  star58_on = 1'b0;
			  star59_on = 1'b0;
			  star60_on = 1'b0;
			  star61_on = 1'b0;
			  star62_on = 1'b0;
			  star63_on = 1'b0;
			  star64_on = 1'b0;
			  star65_on = 1'b0;
			  star66_on = 1'b0;
			  star67_on = 1'b0;
			  star68_on = 1'b0;
			  star69_on = 1'b0;
			  star70_on = 1'b0;
			  star71_on = 1'b0;
			  star72_on = 1'b0;
			  star73_on = 1'b0;
			  star74_on = 1'b0;
			  star75_on = 1'b0;
			  star76_on = 1'b0;
			  star77_on = 1'b0;
			  star78_on = 1'b0;
			  star79_on = 1'b0;
			  star80_on = 1'b0;
			  star81_on = 1'b0;
			  star82_on = 1'b0;
			  star83_on = 1'b0;
			  star84_on = 1'b0;
			  star85_on = 1'b0;
			  star86_on = 1'b0;
			  star87_on = 1'b0;
			  star88_on = 1'b0;
			  star89_on = 1'b0;
			  star90_on = 1'b0;
			  star91_on = 1'b0;
			  star92_on = 1'b0;
			  star93_on = 1'b0;
			  star94_on = 1'b0;
			  star95_on = 1'b0;
			  star96_on = 1'b0;
			  star97_on = 1'b0;
			  star98_on = 1'b0;
			  star99_on = 1'b0;
			  star100_on = 1'b0;
			  star101_on = 1'b0;
			  star102_on = 1'b0;
			  star103_on = 1'b0;
			  star104_on = 1'b0;
			  star105_on = 1'b0;
			  star106_on = 1'b0;
			  star107_on = 1'b0;
			  star108_on = 1'b0;
			  star109_on = 1'b0;
			  star110_on = 1'b0;
			  star111_on = 1'b0;
			  star112_on = 1'b0;
			  star113_on = 1'b0;
			  star114_on = 1'b0;
			  star115_on = 1'b0;
			  star116_on = 1'b0;
			  star117_on = 1'b0;
			  star118_on = 1'b0;
			  star119_on = 1'b0;
			  star120_on = 1'b0;			  
			  ship_addr = (DistY*40 + DistX);
			  alien_addr = 19'b0;
		end
		
		//star 1
	   else if ( ( DistStar1X*DistStar1X + DistStar1Y*DistStar1Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
		   am1_on = 1'b0;
		   am2_on = 1'b0;
		   am3_on = 1'b0;
		   am4_on = 1'b0;
		   am5_on = 1'b0;
		   am6_on = 1'b0;
		   am7_on = 1'b0;
		   am8_on = 1'b0;
		   am9_on = 1'b0;
		   am10_on = 1'b0;
		   am11_on = 1'b0;
		   am12_on = 1'b0;
			star1_on = 1'b1;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;	
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;	
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;	
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 2
	   else if ( ( DistStar2X*DistStar2X + DistStar2Y*DistStar2Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b1;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;	
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 3
	   else if ( ( DistStar3X*DistStar3X + DistStar3Y*DistStar3Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b1;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;	
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;	
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;	
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 4
	   else if ( ( DistStar4X*DistStar4X + DistStar4Y*DistStar4Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b1;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;	
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 5
	   else if ( ( DistStar5X*DistStar5X + DistStar5Y*DistStar5Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
		   am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b1;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;		
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;	
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 6
	   else if ( ( DistStar6X*DistStar6X + DistStar6Y*DistStar6Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b1;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 7
	   else if ( ( DistStar7X*DistStar7X + DistStar7Y*DistStar7Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b1;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;	
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 8
	   else if ( ( DistStar8X*DistStar8X + DistStar8Y*DistStar8Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b1;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 9
	   else if ( ( DistStar9X*DistStar9X + DistStar9Y*DistStar9Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b1;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 10
	   else if ( ( DistStar10X*DistStar10X + DistStar10Y*DistStar10Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b1;
			star11_on = 1'b0;
			star12_on = 1'b0;	
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 11
	   else if ( ( DistStar11X*DistStar11X + DistStar11Y*DistStar11Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b1;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 12
	   else if ( ( DistStar12X*DistStar12X + DistStar12Y*DistStar12Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b1;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;						
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 13
	   else if ( ( DistStar13X*DistStar13X + DistStar13Y*DistStar13Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b1;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 14
	   else if ( ( DistStar14X*DistStar14X + DistStar14Y*DistStar14Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b1;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 15
	   else if ( ( DistStar15X*DistStar15X + DistStar15Y*DistStar15Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b1;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 16
	   else if ( ( DistStar16X*DistStar16X + DistStar16Y*DistStar16Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b1;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 17
	   else if ( ( DistStar17X*DistStar17X + DistStar17Y*DistStar17Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b1;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 18
	   else if ( ( DistStar18X*DistStar18X + DistStar18Y*DistStar18Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b1;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 19
	   else if ( ( DistStar19X*DistStar19X + DistStar19Y*DistStar19Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b1;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 20
	   else if ( ( DistStar20X*DistStar20X + DistStar20Y*DistStar20Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b1;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 21
	   else if ( ( DistStar21X*DistStar21X + DistStar21Y*DistStar21Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b1;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 22
	   else if ( ( DistStar22X*DistStar22X + DistStar22Y*DistStar22Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b1;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 23
	   else if ( ( DistStar23X*DistStar23X + DistStar23Y*DistStar23Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b1;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 24
	   else if ( ( DistStar24X*DistStar24X + DistStar24Y*DistStar24Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b1;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 25
	   else if ( ( DistStar25X*DistStar25X + DistStar25Y*DistStar25Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b1;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 26
	   else if ( ( DistStar26X*DistStar26X + DistStar26Y*DistStar26Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b1;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 27
	   else if ( ( DistStar27X*DistStar27X + DistStar27Y*DistStar27Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b1;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 28
	   else if ( ( DistStar28X*DistStar28X + DistStar28Y*DistStar28Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b1;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 29
	   else if ( ( DistStar29X*DistStar29X + DistStar29Y*DistStar29Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b1;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 30
	   else if ( ( DistStar30X*DistStar30X + DistStar30Y*DistStar30Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b1;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 31
	   else if ( ( DistStar31X*DistStar31X + DistStar31Y*DistStar31Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b1;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 32
	   else if ( ( DistStar32X*DistStar32X + DistStar32Y*DistStar32Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b1;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end	

		//star 33
	   else if ( ( DistStar33X*DistStar33X + DistStar33Y*DistStar33Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b1;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 33
	   else if ( ( DistStar34X*DistStar34X + DistStar34Y*DistStar34Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b1;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 35
	   else if ( ( DistStar35X*DistStar35X + DistStar35Y*DistStar35Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b1;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 36
	   else if ( ( DistStar36X*DistStar36X + DistStar36Y*DistStar36Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b1;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 37
	   else if ( ( DistStar37X*DistStar37X + DistStar37Y*DistStar37Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b1;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 38
	   else if ( ( DistStar38X*DistStar38X + DistStar38Y*DistStar38Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b1;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 39
	   else if ( ( DistStar39X*DistStar39X + DistStar39Y*DistStar39Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b1;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 40
	   else if ( ( DistStar40X*DistStar40X + DistStar40Y*DistStar40Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b1;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 41
	   else if ( ( DistStar41X*DistStar41X + DistStar41Y*DistStar41Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b1;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 42
	   else if ( ( DistStar42X*DistStar42X + DistStar42Y*DistStar42Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b1;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 43
	   else if ( ( DistStar43X*DistStar43X + DistStar43Y*DistStar43Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b1;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 44
	   else if ( ( DistStar44X*DistStar44X + DistStar44Y*DistStar44Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b1;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 45
	   else if ( ( DistStar45X*DistStar45X + DistStar45Y*DistStar45Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b1;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 46
	   else if ( ( DistStar46X*DistStar46X + DistStar46Y*DistStar46Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b1;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 47
	   else if ( ( DistStar47X*DistStar47X + DistStar47Y*DistStar47Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b1;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 48
	   else if ( ( DistStar48X*DistStar48X + DistStar48Y*DistStar48Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b1;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 49
	   else if ( ( DistStar49X*DistStar49X + DistStar49Y*DistStar49Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b1;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 50
	   else if ( ( DistStar50X*DistStar50X + DistStar50Y*DistStar50Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b1;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 51
	   else if ( ( DistStar51X*DistStar51X + DistStar51Y*DistStar51Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b1;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 52
	   else if ( ( DistStar52X*DistStar52X + DistStar52Y*DistStar52Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b1;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 53
	   else if ( ( DistStar53X*DistStar53X + DistStar53Y*DistStar53Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b1;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 54
	   else if ( ( DistStar54X*DistStar54X + DistStar54Y*DistStar54Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b1;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 55
	   else if ( ( DistStar55X*DistStar55X + DistStar55Y*DistStar55Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b1;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 56
	   else if ( ( DistStar56X*DistStar56X + DistStar56Y*DistStar56Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b1;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 57
	   else if ( ( DistStar57X*DistStar57X + DistStar57Y*DistStar57Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b1;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 58
	   else if ( ( DistStar58X*DistStar58X + DistStar58Y*DistStar58Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b1;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 59
	   else if ( ( DistStar59X*DistStar59X + DistStar59Y*DistStar59Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b1;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 60
	   else if ( ( DistStar60X*DistStar60X + DistStar60Y*DistStar60Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b1;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 61
	   else if ( ( DistStar61X*DistStar61X + DistStar61Y*DistStar61Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b1;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 62
	   else if ( ( DistStar62X*DistStar62X + DistStar62Y*DistStar62Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b1;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 63
	   else if ( ( DistStar63X*DistStar63X + DistStar63Y*DistStar63Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b1;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 64
	   else if ( ( DistStar64X*DistStar64X + DistStar64Y*DistStar64Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b1;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 65
	   else if ( ( DistStar65X*DistStar65X + DistStar65Y*DistStar65Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b1;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 66
	   else if ( ( DistStar66X*DistStar66X + DistStar66Y*DistStar66Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b1;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 67
	   else if ( ( DistStar67X*DistStar67X + DistStar67Y*DistStar67Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b1;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 68
	   else if ( ( DistStar68X*DistStar68X + DistStar68Y*DistStar68Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b1;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 69
	   else if ( ( DistStar69X*DistStar69X + DistStar69Y*DistStar69Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b1;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 70
	   else if ( ( DistStar70X*DistStar70X + DistStar70Y*DistStar70Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b1;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 71
	   else if ( ( DistStar71X*DistStar71X + DistStar71Y*DistStar71Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b1;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 72
	   else if ( ( DistStar72X*DistStar72X + DistStar72Y*DistStar72Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b1;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 73
	   else if ( ( DistStar73X*DistStar73X + DistStar73Y*DistStar73Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b1;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 74
	   else if ( ( DistStar74X*DistStar74X + DistStar74Y*DistStar74Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b1;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 75
	   else if ( ( DistStar75X*DistStar75X + DistStar75Y*DistStar75Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b1;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 76
	   else if ( ( DistStar76X*DistStar76X + DistStar76Y*DistStar76Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b1;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 77
	   else if ( ( DistStar77X*DistStar77X + DistStar77Y*DistStar77Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b1;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 78
	   else if ( ( DistStar78X*DistStar78X + DistStar78Y*DistStar78Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b1;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 79
	   else if ( ( DistStar79X*DistStar79X + DistStar79Y*DistStar79Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b1;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 80
	   else if ( ( DistStar80X*DistStar80X + DistStar80Y*DistStar80Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b1;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 81
	   else if ( ( DistStar81X*DistStar81X + DistStar81Y*DistStar81Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b1;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 82
	   else if ( ( DistStar82X*DistStar82X + DistStar82Y*DistStar82Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b1;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 83
	   else if ( ( DistStar83X*DistStar83X + DistStar83Y*DistStar83Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b1;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 84
	   else if ( ( DistStar84X*DistStar84X + DistStar84Y*DistStar84Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b1;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 85
	   else if ( ( DistStar85X*DistStar85X + DistStar85Y*DistStar85Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b1;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 86
	   else if ( ( DistStar86X*DistStar86X + DistStar86Y*DistStar86Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b1;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 87
	   else if ( ( DistStar87X*DistStar87X + DistStar87Y*DistStar87Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b1;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 88
	   else if ( ( DistStar88X*DistStar88X + DistStar88Y*DistStar88Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b1;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 89
	   else if ( ( DistStar89X*DistStar89X + DistStar89Y*DistStar89Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b1;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 90
	   else if ( ( DistStar90X*DistStar90X + DistStar90Y*DistStar90Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b1;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 91
	   else if ( ( DistStar91X*DistStar91X + DistStar91Y*DistStar91Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b1;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 92
	   else if ( ( DistStar92X*DistStar92X + DistStar92Y*DistStar92Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b1;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 93
	   else if ( ( DistStar93X*DistStar93X + DistStar93Y*DistStar93Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b1;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 94
	   else if ( ( DistStar94X*DistStar94X + DistStar94Y*DistStar94Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b1;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 95
	   else if ( ( DistStar95X*DistStar95X + DistStar95Y*DistStar95Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b1;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 96
	   else if ( ( DistStar96X*DistStar96X + DistStar96Y*DistStar96Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b1;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end

		//star 97
	   else if ( ( DistStar97X*DistStar97X + DistStar97Y*DistStar97Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b1;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 98
	   else if ( ( DistStar98X*DistStar98X + DistStar98Y*DistStar98Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b1;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 99
	   else if ( ( DistStar99X*DistStar99X + DistStar99Y*DistStar99Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b1;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 100
	   else if ( ( DistStar100X*DistStar100X + DistStar100Y*DistStar100Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b1;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 101
	   else if ( ( DistStar101X*DistStar101X + DistStar101Y*DistStar101Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b1;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 102
	   else if ( ( DistStar102X*DistStar102X + DistStar102Y*DistStar102Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b1;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 103
	   else if ( ( DistStar103X*DistStar103X + DistStar103Y*DistStar103Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b1;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 104
	   else if ( ( DistStar104X*DistStar104X + DistStar104Y*DistStar104Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b1;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 105
	   else if ( ( DistStar105X*DistStar105X + DistStar105Y*DistStar105Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b1;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 106
	   else if ( ( DistStar106X*DistStar106X + DistStar106Y*DistStar106Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b1;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 107
	   else if ( ( DistStar107X*DistStar107X + DistStar107Y*DistStar107Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b1;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 108
	   else if ( ( DistStar108X*DistStar108X + DistStar108Y*DistStar108Y) <= (star_size * star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b1;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b1;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 109
	   else if ( ( DistStar109X*DistStar109X + DistStar109Y*DistStar109Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b1;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 110
	   else if ( ( DistStar110X*DistStar110X + DistStar110Y*DistStar110Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b1;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 111
	   else if ( ( DistStar111X*DistStar111X + DistStar111Y*DistStar111Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b1;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 112
	   else if ( ( DistStar112X*DistStar112X + DistStar112Y*DistStar112Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b1;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 113
	   else if ( ( DistStar113X*DistStar113X + DistStar113Y*DistStar113Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b1;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 114
	   else if ( ( DistStar114X*DistStar114X + DistStar114Y*DistStar114Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b1;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 115
	   else if ( ( DistStar115X*DistStar115X + DistStar115Y*DistStar115Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b1;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 116
	   else if ( ( DistStar116X*DistStar116X + DistStar116Y*DistStar116Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b1;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 117
	   else if ( ( DistStar117X*DistStar117X + DistStar117Y*DistStar117Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b1;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 118
	   else if ( ( DistStar118X*DistStar118X + DistStar118Y*DistStar118Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b1;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 119
	   else if ( ( DistStar119X*DistStar119X + DistStar119Y*DistStar119Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b1;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//star 120
	   else if ( ( DistStar120X*DistStar120X + DistStar120Y*DistStar120Y) <= (small_star_size * small_star_size) ) 
      begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;	
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b1;		
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
		
		//Alien One
		else if(DrawX >= Alien1X && DrawX < Alien1X + Alien1S &&
			DrawY >= Alien1Y && DrawY < Alien1Y + Alien1S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b1;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;		
			ship_addr = 19'b0;
			alien_addr = (DistAlien1Y*25 + DistAlien1X);
			sprite_addr = 10'b0;
		end
		
		else if(DrawX >= Alien2X && DrawX < Alien2X + Alien2S &&
				DrawY >= Alien2Y && DrawY < Alien2Y + Alien2S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b1;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;			
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;			
			ship_addr = 19'b0;
			alien_addr = (DistAlien2Y*25 + DistAlien2X);
			sprite_addr = 10'b0;
		end
		
		else if(DrawX >= Alien3X && DrawX < Alien3X + Alien3S &&
				DrawY >= Alien3Y && DrawY < Alien3Y + Alien3S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b1;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = (DistAlien3Y*25 + DistAlien3X);			
			sprite_addr = 10'b0;
		end

		else if(DrawX >= Alien4X && DrawX < Alien4X + Alien4S &&
				DrawY >= Alien4Y && DrawY < Alien4Y + Alien4S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b1;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = (DistAlien4Y*25 + DistAlien4X);		
			sprite_addr = 10'b0;
		end

		else if(DrawX >= Alien5X && DrawX < Alien5X + Alien5S &&
				DrawY >= Alien5Y && DrawY < Alien5Y + Alien5S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b1;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = (DistAlien5Y*25 + DistAlien5X);		
			sprite_addr = 10'b0;
		end

		else if(DrawX >= Alien6X && DrawX < Alien6X + Alien6S &&
				DrawY >= Alien6Y && DrawY < Alien6Y + Alien6S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b1;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = (DistAlien6Y*25 + DistAlien6X);		
			sprite_addr = 10'b0;
		end
		
		else if(DrawX >= Alien7X && DrawX < Alien7X + Alien7S &&
				DrawY >= Alien7Y && DrawY < Alien7Y + Alien7S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b1;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = (DistAlien7Y*25 + DistAlien7X);		
			sprite_addr = 10'b0;
		end
		
		else if(DrawX >= Alien8X && DrawX < Alien8X + Alien8S &&
				DrawY >= Alien8Y && DrawY < Alien8Y + Alien8S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b1;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			ship_addr = 19'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			alien_addr = (DistAlien8Y*25 + DistAlien8X);		
			sprite_addr = 10'b0;
		end	
		
		else if(DrawX >= Alien9X && DrawX < Alien9X + Alien9S &&
				DrawY >= Alien9Y && DrawY < Alien9Y + Alien9S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b1;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			ship_addr = 19'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			alien_addr = (DistAlien9Y*25 + DistAlien9X);		
			sprite_addr = 10'b0;
		end
	
		else if(DrawX >= Alien10X && DrawX < Alien10X + Alien10S &&
				DrawY >= Alien10Y && DrawY < Alien10Y + Alien10S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b1;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			ship_addr = 19'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			alien_addr = (DistAlien10Y*25 + DistAlien10X);		
			sprite_addr = 10'b0;
		end
	
		else if(DrawX >= Alien11X && DrawX < Alien11X + Alien11S &&
				DrawY >= Alien11Y && DrawY < Alien11Y + Alien11S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b1;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = (DistAlien11Y*25 + DistAlien11X);		
			sprite_addr = 10'b0;
		end

		else if(DrawX >= Alien12X && DrawX < Alien12X + Alien12S &&
				DrawY >= Alien12Y && DrawY < Alien12Y + Alien12S)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b1;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = (DistAlien12Y*25 + DistAlien12X);		
			sprite_addr = 10'b0;
		end
		
		else if(DrawX >= MissileX && DrawX < MissileX + MissileS &&
				DrawY >= MissileY && DrawY < MissileY + 2*MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b1;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end
		
		//Draw AM1
		else if(DrawX >= Alien1MissileX && DrawX < Alien1MissileX + Alien1MissileS &&
				DrawY >= Alien1MissileY && DrawY < Alien1MissileY + 2*Alien1MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b1;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM2
		else if(DrawX >= Alien2MissileX && DrawX < Alien2MissileX + Alien2MissileS &&
				DrawY >= Alien2MissileY && DrawY < Alien2MissileY + 2*Alien2MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b1;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM3
		else if(DrawX >= Alien3MissileX && DrawX < Alien3MissileX + Alien3MissileS &&
				DrawY >= Alien3MissileY && DrawY < Alien3MissileY + 2*Alien3MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b1;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM4
		else if(DrawX >= Alien4MissileX && DrawX < Alien4MissileX + Alien4MissileS &&
				DrawY >= Alien4MissileY && DrawY < Alien4MissileY + 2*Alien4MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b1;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM5
		else if(DrawX >= Alien5MissileX && DrawX < Alien5MissileX + Alien5MissileS &&
				DrawY >= Alien5MissileY && DrawY < Alien5MissileY + 2*Alien5MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b1;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM6
		else if(DrawX >= Alien6MissileX && DrawX < Alien6MissileX + Alien6MissileS &&
				DrawY >= Alien6MissileY && DrawY < Alien6MissileY + 2*Alien6MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b1;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM7
		else if(DrawX >= Alien7MissileX && DrawX < Alien7MissileX + Alien7MissileS &&
				DrawY >= Alien7MissileY && DrawY < Alien7MissileY + 2*Alien7MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b1;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM1
		else if(DrawX >= Alien8MissileX && DrawX < Alien8MissileX + Alien8MissileS &&
				DrawY >= Alien8MissileY && DrawY < Alien8MissileY + 2*Alien8MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b1;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM9
		else if(DrawX >= Alien9MissileX && DrawX < Alien9MissileX + Alien9MissileS &&
				DrawY >= Alien9MissileY && DrawY < Alien9MissileY + 2*Alien9MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b1;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM10
		else if(DrawX >= Alien10MissileX && DrawX < Alien10MissileX + Alien10MissileS &&
				DrawY >= Alien10MissileY && DrawY < Alien10MissileY + 2*Alien10MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b1;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM11
		else if(DrawX >= Alien11MissileX && DrawX < Alien11MissileX + Alien11MissileS &&
				DrawY >= Alien11MissileY && DrawY < Alien11MissileY + 2*Alien11MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b1;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Draw AM12
		else if(DrawX >= Alien12MissileX && DrawX < Alien12MissileX + Alien12MissileS &&
				DrawY >= Alien12MissileY && DrawY < Alien12MissileY + 2*Alien12MissileS)
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b1;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;;
		end

		//Default Zero Value 
		else
		begin
			ball_on = 1'b0;
			alien1_on = 1'b0;
			alien2_on = 1'b0;
			alien3_on = 1'b0;
			alien4_on = 1'b0;
			alien5_on = 1'b0;
			alien6_on = 1'b0;
			alien7_on = 1'b0;
		   alien8_on = 1'b0;
		   alien9_on = 1'b0;
		   alien10_on = 1'b0;
		   alien11_on = 1'b0;
		   alien12_on = 1'b0;
			missile_on = 1'b0;
			am1_on = 1'b0;
			am2_on = 1'b0;
			am3_on = 1'b0;
			am4_on = 1'b0;
			am5_on = 1'b0;
			am6_on = 1'b0;
			am7_on = 1'b0;
			am8_on = 1'b0;
		   am9_on = 1'b0;
			am10_on = 1'b0;
			am11_on = 1'b0;
			am12_on = 1'b0;
			star1_on = 1'b0;
			star2_on = 1'b0;
			star3_on = 1'b0;
			star4_on = 1'b0;
			star5_on = 1'b0;
			star6_on = 1'b0;
			star7_on = 1'b0;
			star8_on = 1'b0;
			star9_on = 1'b0;
			star10_on = 1'b0;
			star11_on = 1'b0;
			star12_on = 1'b0;
			star13_on = 1'b0;
			star14_on = 1'b0;
			star15_on = 1'b0;
			star16_on = 1'b0;
			star17_on = 1'b0;
			star18_on = 1'b0;
			star19_on = 1'b0;
			star20_on = 1'b0;
			star21_on = 1'b0;
			star22_on = 1'b0;
			star23_on = 1'b0;
			star24_on = 1'b0;
			star25_on = 1'b0;
			star26_on = 1'b0;
			star27_on = 1'b0;
			star28_on = 1'b0;
			star29_on = 1'b0;
			star30_on = 1'b0;
			star31_on = 1'b0;
			star32_on = 1'b0;
			star33_on = 1'b0;
			star34_on = 1'b0;
			star35_on = 1'b0;
			star36_on = 1'b0;
			star37_on = 1'b0;
			star38_on = 1'b0;
			star39_on = 1'b0;
			star40_on = 1'b0;
			star41_on = 1'b0;
			star42_on = 1'b0;
			star43_on = 1'b0;
			star44_on = 1'b0;
			star45_on = 1'b0;
			star46_on = 1'b0;
			star47_on = 1'b0;
			star48_on = 1'b0;
			star49_on = 1'b0;
			star50_on = 1'b0;
			star51_on = 1'b0;
			star52_on = 1'b0;
			star53_on = 1'b0;
			star54_on = 1'b0;
			star55_on = 1'b0;
			star56_on = 1'b0;
			star57_on = 1'b0;
			star58_on = 1'b0;
			star59_on = 1'b0;
			star60_on = 1'b0;
			star61_on = 1'b0;
			star62_on = 1'b0;
			star63_on = 1'b0;
			star64_on = 1'b0;
			star65_on = 1'b0;
			star66_on = 1'b0;
			star67_on = 1'b0;
			star68_on = 1'b0;
			star69_on = 1'b0;
			star70_on = 1'b0;
			star71_on = 1'b0;
			star72_on = 1'b0;
			star73_on = 1'b0;
			star74_on = 1'b0;
			star75_on = 1'b0;
			star76_on = 1'b0;
			star77_on = 1'b0;
			star78_on = 1'b0;
			star79_on = 1'b0;
			star80_on = 1'b0;
			star81_on = 1'b0;
			star82_on = 1'b0;
			star83_on = 1'b0;
			star84_on = 1'b0;
			star85_on = 1'b0;
			star86_on = 1'b0;
			star87_on = 1'b0;
			star88_on = 1'b0;
			star89_on = 1'b0;
			star90_on = 1'b0;
			star91_on = 1'b0;
			star92_on = 1'b0;
			star93_on = 1'b0;
			star94_on = 1'b0;
			star95_on = 1'b0;
			star96_on = 1'b0;
			star97_on = 1'b0;
			star98_on = 1'b0;
			star99_on = 1'b0;
			star100_on = 1'b0;
			star101_on = 1'b0;
			star102_on = 1'b0;
			star103_on = 1'b0;
			star104_on = 1'b0;
			star105_on = 1'b0;
			star106_on = 1'b0;
			star107_on = 1'b0;
			star108_on = 1'b0;
			star109_on = 1'b0;
			star110_on = 1'b0;
			star111_on = 1'b0;
			star112_on = 1'b0;
			star113_on = 1'b0;
			star114_on = 1'b0;
			star115_on = 1'b0;
			star116_on = 1'b0;
			star117_on = 1'b0;
			star118_on = 1'b0;
			star119_on = 1'b0;
			star120_on = 1'b0;
			ship_addr = 19'b0;
			alien_addr = 19'b0;		
			sprite_addr = 10'b0;
		end
	 end 
	 
    always_comb
    begin:RGB_Display
	     if ((ball_on == 1'b1)) 
        begin 
            Red = dout[23:16];
            Green = dout[15:8];            
			   Blue = dout[7:0];
        end 
		  
        else if ((alien1_on == 1'b1) && (alien1_hit == 0)) 
        begin 
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
        end  
		  
		  else if((alien2_on == 1'b1) && (alien2_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end

		  else if((alien3_on == 1'b1) && (alien3_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end
		  
		  else if((alien4_on == 1'b1) && (alien4_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];		  
		  end
		  
		  else if((alien5_on == 1'b1) && (alien5_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end
		  
		  else if((alien6_on == 1'b1) && (alien6_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end

		  else if((alien7_on == 1'b1) && (alien7_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end
		  
		  else if((alien8_on == 1'b1) && (alien8_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end
		  
		  else if((alien9_on == 1'b1) && (alien9_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end
		  
		  else if((alien10_on == 1'b1) && (alien10_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end
		  
		  else if((alien11_on == 1'b1) && (alien11_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end
		   
		  else if((alien12_on == 1'b1) && (alien12_hit == 0))
		  begin
            Red = dout_1[23:16];
            Green = dout_1[15:8];            
			   Blue = dout_1[7:0];
		  end
		  
		  else if((missile_on == 1'b1) && (missile_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'hff;
            Blue = 8'h00;
		  end
		  
		  else if((am1_on == 1'b1) && (am1_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am2_on == 1'b1) && (am2_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am3_on == 1'b1) && (am3_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am4_on == 1'b1) && (am4_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am5_on == 1'b1) && (am5_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am6_on == 1'b1) && (am6_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am7_on == 1'b1) && (am7_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am8_on == 1'b1) && (am8_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am9_on == 1'b1) && (am9_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am10_on == 1'b1) && (am10_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am11_on == 1'b1) && (am11_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((am12_on == 1'b1) && (am12_sight == 1'b1))
		  begin
            Red = 8'hff;
            Green = 8'h80;
            Blue = 8'h00;
		  end
		  
		  else if((star1_on == 1'b1) || (star2_on == 1'b1) || (star3_on == 1'b1) || (star4_on == 1'b1) || (star5_on == 1'b1)
						|| (star6_on == 1'b1) || (star7_on == 1'b1) || (star8_on == 1'b1) || (star9_on == 1'b1) || (star10_on == 1'b1) || (star11_on == 1'b1) || (star12_on == 1'b1)
						|| (star25_on == 1'b1) || (star26_on == 1'b1) || (star27_on == 1'b1) || (star28_on == 1'b1) || (star29_on == 1'b1) || (star30_on == 1'b1) || (star31_on == 1'b1)
						|| (star32_on == 1'b1) || (star33_on == 1'b1) || (star34_on == 1'b1) || (star35_on == 1'b1) || (star36_on == 1'b1)
						|| (star49_on == 1'b1) || (star50_on == 1'b1) || (star51_on == 1'b1) || (star52_on == 1'b1) || (star53_on == 1'b1) || (star54_on == 1'b1) || (star55_on == 1'b1)
						|| (star56_on == 1'b1) || (star57_on == 1'b1) || (star58_on == 1'b1) || (star59_on == 1'b1) || (star60_on == 1'b1)
						|| (star73_on == 1'b1) || (star74_on == 1'b1) || (star75_on == 1'b1) || (star76_on == 1'b1) || (star77_on == 1'b1) || (star78_on == 1'b1) || (star79_on == 1'b1)
						|| (star80_on == 1'b1) || (star81_on == 1'b1) || (star82_on == 1'b1) || (star83_on == 1'b1) || (star84_on == 1'b1)
						|| (star97_on == 1'b1) || (star98_on == 1'b1) || (star99_on == 1'b1) || (star100_on == 1'b1) || (star101_on == 1'b1) || (star102_on == 1'b1) || (star103_on == 1'b1)
						|| (star104_on == 1'b1) || (star105_on == 1'b1) || (star106_on == 1'b1) || (star107_on == 1'b1) || (star108_on == 1'b1))
		  begin
				if(color_switch)
				begin
					Red = 8'hff;
					Green = 8'h00;
					Blue = 8'h00;
				end
				else
				begin
					Red = 8'he0;
					Green = 8'he0;
					Blue = 8'he0;
				end
		  end
		  
		  else if((star13_on == 1'b1) || (star14_on == 1'b1) || (star15_on == 1'b1) || (star16_on == 1'b1) || (star17_on == 1'b1)
						|| (star18_on == 1'b1) || (star19_on == 1'b1) || (star20_on == 1'b1) || (star21_on == 1'b1) || (star22_on == 1'b1) || (star23_on == 1'b1) || (star24_on == 1'b1)
						|| (star37_on == 1'b1) || (star38_on == 1'b1) || (star39_on == 1'b1) || (star40_on == 1'b1) || (star41_on == 1'b1) || (star42_on == 1'b1) || (star43_on == 1'b1)
						|| (star44_on == 1'b1) || (star45_on == 1'b1) || (star46_on == 1'b1) || (star47_on == 1'b1) || (star48_on == 1'b1)
						|| (star61_on == 1'b1) || (star62_on == 1'b1) || (star63_on == 1'b1) || (star64_on == 1'b1) || (star65_on == 1'b1) || (star66_on == 1'b1) || (star67_on == 1'b1)
						|| (star68_on == 1'b1) || (star69_on == 1'b1) || (star70_on == 1'b1) || (star71_on == 1'b1) || (star72_on == 1'b1)
						|| (star85_on == 1'b1) || (star86_on == 1'b1) || (star87_on == 1'b1) || (star88_on == 1'b1) || (star89_on == 1'b1) || (star90_on == 1'b1) || (star91_on == 1'b1)
						|| (star92_on == 1'b1) || (star93_on == 1'b1) || (star94_on == 1'b1) || (star95_on == 1'b1) || (star96_on == 1'b1)
						|| (star109_on == 1'b1) || (star110_on == 1'b1) || (star111_on == 1'b1) || (star112_on == 1'b1) || (star113_on == 1'b1) || (star114_on == 1'b1) || (star115_on == 1'b1)
						|| (star116_on == 1'b1) || (star117_on == 1'b1) || (star118_on == 1'b1) || (star119_on == 1'b1) || (star120_on == 1'b1))
		  begin
			if(color_switch)
				begin
					Red = 8'h00;
					Green = 8'h80;
					Blue = 8'hff;
				end
				else
				begin
					Red = 8'he0;
					Green = 8'he0;
					Blue = 8'he0;
				end
		  end
		  
        else  
        begin 
            Red = 8'h00; 
            Green = 8'h00;
            Blue = 8'h00;
       end      
    end 
	 
endmodule
